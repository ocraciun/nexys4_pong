library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity driver7seg is
    Port ( CLK : in STD_LOGIC; --100MHz board clock input
           Din : in STD_LOGIC_VECTOR (31 downto 0); --31 bit binary data for 4 displays
           an : out STD_LOGIC_VECTOR (7 downto 0); --anode outputs selecting individual displays 7 to 0
           seg : out STD_LOGIC_VECTOR (0 to 6); -- cathode outputs for selecting LED-s in each display
           dp_in : in STD_LOGIC_VECTOR (7 downto 0); --decimal point input values
           dp_out : out STD_LOGIC; --selected decimal point sent to cathodes
           RST : in STD_LOGIC); --global reset
end driver7seg;

architecture Behavioral of driver7seg is

signal clk1kHz : STD_LOGIC;
signal state : STD_LOGIC_VECTOR(16 downto 0);
signal addr : STD_LOGIC_VECTOR(2 downto 0);
signal cseg : STD_LOGIC_VECTOR(3 downto 0);

begin

-- frequency divider by 100k to generate 1kHz anode sweeping clock
-- counting from 0 to 99999, output is MSB 
-- 17 counter state length needed 
div1kHz: process(CLK, RST)
begin
   if RST = '0' then 
        state <= '0' & X"0000";
   else
     if rising_edge(CLK) then
        if state = '1' & X"869F" then --if counte reaches 99999
            state <= '0' & X"0000"; -- reset back to 0
        else
            state <= state+1;
        end if;
     end if;
   end if;         
end process;

clk1Khz <= state(16); --assign MSB to frequency divider output


-- 2 bit counter generating 4 addresses for display multiplexing
counter_2bits: process(clk1kHz)
begin
  if rising_edge(clk1kHz) then       
           addr <= addr+1;   
  end if;   
end process;

-- 3 to 8 decoder used to select one display of 8 at each sweeping address generated by the 3 bit counter 
-- anodes are active low, decoder must provide '0' for activation
dcd3_8: process(addr)
begin
  case addr is
      when "000" =>  an <= "01111111";       
      when "001" =>  an <= "10111111"; 
      when "010" =>  an <= "11011111"; 
      when "011" =>  an <= "11101111";
      when "100" =>  an <= "11110111";       
      when "101" =>  an <= "11111011"; 
      when "110" =>  an <= "11111101"; 
      when "111" =>  an <= "11111110";  
      when others => an <= "11111111";
   end case; 
end process;

--4 input multiplexer to select data to be sent to a single display
--synchronzied with addr and display activation with the anodes
data_mux4: process(addr,Din,dp_in)
begin
  case addr is
      when "000" =>  cseg <= Din(31 downto 28); -- sending 4 upper bits targeted at display 7 
                    dp_out <= not dp_in(7);     -- lighting up decimal point on display 7
      when "001" =>  cseg <= Din(27 downto 24); -- sending next 4 bits targeted at display 6
                    dp_out <= not dp_in(6);     -- lighting up decimal point on display 6
      when "010" =>  cseg <= Din(23 downto 20); -- sending 4 upper bits targeted at display 5 
                    dp_out <= not dp_in(5);     -- lighting up decimal point on display 5
      when "011" =>  cseg <= Din(19 downto 16); -- sending 4 upper bits targeted at display 4 
                    dp_out <= not dp_in(4);     -- lighting up decimal point on display 4
      when "100" =>  cseg <= Din(15 downto 12); -- sending 4 upper bits targeted at display 3  
                    dp_out <= not dp_in(3);     -- lighting up decimal point on display 3
      when "101" =>  cseg <= Din(11 downto 8);  -- sending next 4 bits targeted at display 2
                    dp_out <= not dp_in(2);     -- lighting up decimal point on display 2
      when "110" =>  cseg <= Din(7 downto 4);   -- sending 4 upper bits targeted at display 1 
                    dp_out <= not dp_in(1);     -- lighting up decimal point on display 1
      when "111" =>  cseg <= Din(3 downto 0);   -- sending 4 upper bits targeted at display 0 
                    dp_out <= not dp_in(0);     -- lighting up decimal point on display 0
      when others => cseg <= "XXXX";
                     dp_out <= 'X';
   end case; 
end process;

--binary to 7 segment decoder
--cathodes also active low, provide '0' for a lit up segment or decimal point
dcd7seg:process(cseg)
begin
  case cseg is
      when "0000" =>  seg <= "0000001"; -- 0
      when "0001" =>  seg <= "1001111"; -- 1
      when "0010" =>  seg <= "0010010"; -- 2
      when "0011" =>  seg <= "0000110"; -- 3
      when "0100" =>  seg <= "1001100"; -- 4
      when "0101" =>  seg <= "0100100"; -- 5
      when "0110" =>  seg <= "0100000"; -- 6
      when "0111" =>  seg <= "0001111"; -- 7
      when "1000" =>  seg <= "0000000"; -- 8
      when "1001" =>  seg <= "0000100"; -- 9
      --when "1010" =>  seg <= "0000010"; -- A
     -- when "1011" =>  seg <= "1100000"; -- B
      --when "1100" =>  seg <= "0110001"; -- C
      --when "1101" =>  seg <= "1000010"; -- D
      --when "1110" =>  seg <= "0110000"; -- E
      --when "1111" =>  seg <= "0111000"; -- F
      when others =>  seg <= "0011000"; -- P
   end case; 
end process;

end Behavioral;
