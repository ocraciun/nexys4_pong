`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/20/2023 07:37:43 PM
// Design Name: 
// Module Name: pong_game
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module pong_game(
    input CLK,
    output [3:0] VGA_RED_O,
    output [3:0] VGA_GREEN_O,
    output [3:0] VGA_BLUE_O,
    output VGA_H_SYNC_O,
    output VGA_V_SYNC_O
    );
endmodule
